module demux (output logic [7:0] Y, input logic D, input logic [2:0] SEL);
  
  
endmodule

